 /*                                                                      
 Copyright 2020 Blue Liang, liangkangnan@163.com
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
 Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */

`include "include.v"


// 32 bits count up timer module
module timer(

    input wire clk,
    input wire rst_n,

    input wire[31:0] data_i,
    input wire[31:0] addr_i,
    input req_i,
    input wire we_i,

    output addr_ok,
    output data_ok,
    input [`RAM_MASK_WIDTH - 1: 0]wem,

    output reg[31:0] data_o,
    output wire int_sig_o

    );

    localparam REG_CTRL = 4'h0;
    localparam REG_COUNT = 4'h4;
    localparam REG_VALUE = 4'h8;

    reg read_data_ok;
    reg write_data_ok;
    assign addr_ok = req_i;
    assign data_ok = read_data_ok | write_data_ok;
    // [0]: timer enable
    // [1]: timer int enable
    // [2]: timer int pending, write 1 to clear it
    // addr offset: 0x00
    reg[31:0] timer_ctrl;

    // timer current count, read only
    // addr offset: 0x04
    reg[31:0] timer_count;

    // timer expired value
    // addr offset: 0x08
    reg[31:0] timer_value;


    assign int_sig_o = ((timer_ctrl[2] == 1'b1) && (timer_ctrl[1] == 1'b1))? `INT_ASSERT: `INT_DEASSERT;

    // counter
	always@(posedge clk )begin
        if (!rst_n) begin
            timer_count <= 0;
        end else begin
            if (timer_ctrl[0] == 1'b1) begin
                timer_count <= timer_count + 1'b1;
                if (timer_count >= timer_value) begin
                    timer_count <=  0;
                end
            end else begin
                timer_count <=  0;
            end
        end
    end

    // write regs
	always@(posedge clk)begin
        if (!rst_n) begin
            timer_ctrl <= 0;
            timer_value <=  0;
            write_data_ok <= 1'b0;
        end else if(req_i)begin
            if (we_i) begin
                write_data_ok <= 1'b1;
                case (addr_i[3:0])
                    REG_CTRL: begin
                        timer_ctrl <= {data_i[31:3], (timer_ctrl[2] & (~data_i[2])), data_i[1:0]};
                    end
                    REG_VALUE: begin
                        timer_value <= data_i;
                    end
                endcase
            end else begin
                if ((timer_ctrl[0] == 1'b1) && (timer_count >= timer_value)) begin
                    timer_ctrl[0] <= 1'b0;
                    timer_ctrl[2] <= 1'b1;
                end
            end
        end
        else begin
            write_data_ok <= 1'b0;
        end
    end

    // read regs
	always@(posedge clk)begin
        if (!rst_n) begin
            data_o <= 0;
            read_data_ok <= 1'b0;
        end else if(addr_ok) begin
            read_data_ok <= 1'b1;
            case (addr_i[3:0])
                REG_VALUE: begin
                    data_o <= timer_value;
                end
                REG_CTRL: begin
                    data_o <= timer_ctrl;
                end
                REG_COUNT: begin
                    data_o <= timer_count;
                end
                default: begin
                    data_o <= 0;
                end
            endcase
        end
    end

endmodule
