
module alucontrol(


);
	

endmodule
