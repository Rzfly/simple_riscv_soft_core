
module control(
	input [`DATA_WIDTH]instruction,
	output write_reg,
	output ALU_src,
	output [`ALU_OP_WIDTH]ALU_op,
	output mem2reg,
	output read_mem,
	output write_mem,

);

	

endmodule