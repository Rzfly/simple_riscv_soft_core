`include "include.v"

module hazard_detection(
);

	
endmodule