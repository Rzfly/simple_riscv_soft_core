

`include "include.v"

module branch_addr_gen(
	input [`DATA_WIDTH - 1:0]pc,
	input [`DATA_WIDTH - 1:0]imm,
	output [`DATA_WIDTH - 1:0]branch_addr
);
	
	assign branch_addr = pc + imm;

endmodule